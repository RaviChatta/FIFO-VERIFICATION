
package fifo_pkg;
	import uvm_pkg::*;
	
	`include "uvm_macros.svh"
       	`include "trans.sv"
	`include "sequence.sv"
	`include "sequencer.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "agent.sv"
	`include "scoreboard.sv"
	`include "env.sv"
	`include "test.sv"

endpackage

